`include "structs.sv"

